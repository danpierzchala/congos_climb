------------------------------
------------------------------
--- TOP LEVEL CONGOS CLIMB ---
------------------------------
------------------------------
-- By: Dan Pierzchala 		--
-- and 						--
-- James Rey				--
------------------------------
------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library work;
use work.array_platPos.all;
--------------------------
-- The top level entity of this game has the basic inputs, clock, reset, ps2clock and ps2data
-- and outputs the typical signals needed to display on VGA, the normal hex driver signals are also used
-- to display the score on the 7 segment hex displays
-------------------------

entity toplevel_jumper is
    Port ( Clk 			: in std_logic; -- 50 MHz system clock
           Reset 		: in std_logic; -- global reset
           Red   		: out std_logic_vector(9 downto 0); -- VGA display
           Green 		: out std_logic_vector(9 downto 0); -- VGA display
           Blue  		: out std_logic_vector(9 downto 0); -- VGA display
           VGA_clk 		: out std_logic; -- VGA display 
           sync 		: out std_logic; -- VGA display
           blank 		: out std_logic; -- VGA display
           vs 			: out std_logic; -- VGA display
           hs 			: out std_logic; -- VGA display
           ps2Clk 		: in std_logic; -- PS2 port
           ps2Data 		: in std_logic; -- PS2 port
		   AhexU 		: out std_logic_vector(6 downto 0); -- 7 segment hex display
		   AhexL 		: out std_logic_vector(6 downto 0); -- 7 segment hex display
		   BhexU 		: out std_logic_vector(6 downto 0); -- 7 segment hex display
		   BhexL 		: out std_logic_vector(6 downto 0)); -- 7 segment hex display          	           
end toplevel_jumper;

architecture Behavioral of toplevel_jumper is

------------------------
-- The vga_display_engine is in charge of displaying the current game state to the screen
-- The engine has the basic clock and reset inputs, as well as some position data inputs and directional data inputs
-- Congos X and Y position, and the X and Y platform positions, and the X and Y banana positions are used to draw them to the screen.
-- Because the platform width is not constant, it must also be used as an input to draw the platforms correctly on the screen
-- The the left direction and right direction are used to display the correct sprite on the screen
--
-- The vga_display engine has the normal outputs necessary for correct VGA display, 
-- and also outputs the frame start when a new frame is drawn
------------------------
component vga_display_engine is 
  Port ( clk       	: in  std_logic;  -- 50 MHz system clock
         reset     	: in  std_logic;  -- global reset
         guyPosX	: in std_logic_vector(9 downto 0); -- Congo's x position
         guyPosY	: in std_logic_vector(9 downto 0); -- Congo's y position
         platXpos	: in platArray; -- array of 8 x platform locations
         platYpos1 	: in platArray; -- first array of 8 y platform locations
         platYpos2	: in platArray; -- second array of 8 y platform locations
         platWidth  : in std_logic_vector(9 downto 0); -- platform width
		leftDir		: in std_logic; -- if Congo's moving left, 1
		rightDir	: in std_logic; -- if Congo's moving right, 1
		banPosX		: in std_logic_vector(9 downto 0);
        banPosY		: in std_logic_vector(9 downto 0);
         
         hs        : out std_logic;  -- Horizontal sync pulse.  Active low
         vs        : out std_logic;  -- Vertical sync pulse.  Active low
         pixel_clk : out std_logic;  -- 25 MHz pixel clock output
         blank     : out std_logic;  -- Blanking interval indicator.  Active low.
         sync      : out std_logic;  -- Composite Sync signal.  Active low.  We don't use it in this lab,
                                     --   but the video DAC on the DE2 board requires an input for it.
         fStart		: out std_logic; -- frame start signal
         Red   		: out std_logic_vector(9 downto 0);
         Green 		: out std_logic_vector(9 downto 0);
         Blue  		: out std_logic_vector(9 downto 0));
end component;

---------------------
-- The physics_engine is where the brain of the game is
-- It has the basic clock and reset inputs, a frame start signal, and 
-- left and right inputs from the Congo entity. The physics engine
-- is to process user input and correctly pilot Congo in the game
-- and update his position accordingly, checking collisions with
-- platforms, and making sure he stays visible in the x range of the screen
-- If Congo falls to the bottom of the screen, the physics_engine is stopped and the game is ended
--
--The engine keeps track internally of the bananas and platform positions, both being generated by
-- a platform_generator and a banana_generator. The physics engine is in charge of outputting those positions
-- to the display engine in order to display them correctly on the screen
--
--The engine also keeps track of bananas hit and platforms hit, and outputs the corresponding points gained from them
-- to be sent to the display engine for correct display on the 7seg hex displays
--------------------
component physics_engine is
    Port ( clk		: in std_logic; -- 50 MHz system clock
           Reset	: in std_logic; -- global reset
           fStart	: in std_logic; -- frame start signal from display_engine
           L		: in std_logic; -- From Congo entity, 1 if A pressed
           R		: in std_logic; -- From Congo entity, 1 if D pressed
      
           platw	: out std_logic_vector(9 downto 0);
           dead		: out std_logic; -- dead signal, 1 if Congo fell to the bottom of the screen
           guyPosX	: out std_logic_vector(9 downto 0); -- Congo's x position
           guyPosY	: out std_logic_vector(9 downto 0); -- Congo's y position
           bananaPosX : out std_logic_vector(9 downto 0); -- x position of the banana
           bananaPosY : out std_logic_vector(9 downto 0); -- y position of the banana
           score	: out std_logic_vector(7 downto 0); -- score gained from bananas
           platPosX	: out platArray; -- array of 8 x platform locations
           platPosY1: out platArray; -- first array of 8 y platform locations
           platPosY2: out platArray; -- second array of 8 y platform locations
           jCount	: out std_logic_vector(7 downto 0)); -- total number of platforms hit
end component;


--------------------
-- The guy engine is where the keyboard gets processed and outputs the correct directional signal
-- based on whether A or D was pressed
-- It runs on the system clock and has the global reset signals, and the necessary input signals from the keyboard entity
--------------------
component guy is	
	Port ( clk	: in std_logic; -- 50 MHz system clock
           Reset	: in std_logic; -- global reset signal
           makeIn   : in std_logic; -- from keyboard when new make signal recieved
           codeRdyIn: in std_logic; -- 0->1 when new signal is recieved
           scanIn	: in std_logic_vector(7 downto 0); -- make code
           L		: out std_logic; -- outputs a 1 if A pressed
           R		: out std_logic); -- outputs a 1 if D pressed
end component;	


-------------------
-- The keyboard processor is in charge of reading the data from the ps2 port
-- and collecting the correct make code when a key is pressed
-- It runs on the system clock and has the global reset signal
-- Outputs the scancode, make, and codeRdy signals to the guy unit
-- in order to create the directional signals
------------------
component keyboard is 
   Port ( 
			Clk 	:		in std_logic; -- 50 MHz global clock
			reset 	: 		in std_logic; -- global reset
           psClk	: 		in std_logic; -- PS2 keyboard clock  
           psData 	: 		in std_logic; -- PS2 keyboard data
		   scanCode :	out std_logic_vector(7 downto 0); -- make code
		   codeRdy: 	out std_logic; -- 0->1 if makecode read
		   make:   out std_logic); -- 1 if make code read
end component;
	
--------------------
-- Used for displaying the score on the 7seg hex displays
--------------------
component HexDriver is 
	port ( In0 : in std_logic_vector(3 downto 0);
		   Out0 : out std_logic_vector(6 downto 0));
end component HexDriver;




signal vsSig, Reset_h, fStartSig : std_logic;
signal DrawXSig, DrawYSig, platXsig, platYsig : std_logic_vector(9 downto 0);
signal redSig, greenSig, blueSig : std_logic_vector(9 downto 0);



signal wPlat, wHalfPlat, xGuy, yGuy, sGuy : std_logic_vector(9 downto 0);
signal makeSig, codeReadySig : std_logic;
signal scanCodeSig : std_logic_vector(7 downto 0);

signal xPlatSig, yPlatSig1, yPlatSig2 : platArray;
signal deadsig : std_logic;
signal moveLeftSig, moveRightSig : std_logic;
signal moveLeftVec, moveRightVec, fStartVec : std_logic_vector(3 downto 0);

signal jCountSig, bCountSig	: std_logic_vector(7 downto 0);
signal scoreSig	: std_logic_vector(15 downto 0);


signal guyPosYsig, guyPosXsig : std_logic_vector(9 downto 0);
signal bananaPosYsig, bananaPosXsig : std_logic_vector(9 downto 0);
signal pWidthSig	: std_logic_vector(9 downto 0);




begin

Reset_h <= not Reset;
fStartVec <= "000" & fStartSig;

scoreSig <= ("00000000" & bCountSig) + ("00000000" & jCountSig);

vga_Sync : vga_display_engine
  Port map ( clk       => clk,
         reset     => Reset_h,
         guyPosX   => guyPosXsig,	
         guyPosY	=>	guyPosYsig,	
         platXpos	=> xPlatSig,
         platYpos1 	=> yPlatSig1,
         platYpos2	=> yPlatSig2,
         platWidth	=> pWidthSig,
		leftDir		=> moveLeftSig,
        rightDir	=> moveRightSig,
        banPosX		=> bananaPosXsig,
         banPosY	=> bananaPosYsig,
        
         
         hs        => hs, 
         vs        => vsSig,
         pixel_clk => VGA_clk,
         blank     => blank,
         sync      => sync,                                 
         fStart		=>	fStartSig,
         Red   		=> redSig,
         Green 		=> greenSig,
         Blue  		=> blueSig);
				
game_physics : physics_engine
    Port Map(clk	=> clk,
           Reset	=> Reset_h,
           fStart	=> fStartSig,
           L		=> moveLeftSig,
           R		=> moveRightSig,
           
           platW	=> pWidthSig,
           score	=> bCountSig,
           dead		=> deadSig,
           guyPosX	=> guyPosXsig, 
           guyPosY	=> guyPosYsig, 
           bananaPosX => bananaPosXsig,
           bananaPosY => bananaPosYsig, 
           platPosX	=> xPlatSig,
           platPosY1=> yPlatSig1,
           platPosY2=> yPlatSig2,
           jCount	=> jCountSig);
				
guy_instance : guy
	Port Map(  clk	=> vsSig,
				Reset	=> Reset_h,
				scanIn => scanCodeSig,
				makeIn => makeSig,
				codeRdyIn => codeReadySig,
				L => moveLeftSig,
				R => moveRightSig);
				
keyboard_instance : keyboard
	Port Map( 	Clk 	=> Clk,
				reset 	=> Reset_h,
			   psClk	=> ps2Clk,	
			   psData 	=> ps2Data,		
			   scanCode => scanCodeSig,
			   codeRdy => codeReadySig,
			   make     => makeSig);
			   
HexA_U : HexDriver
	port map ( In0 => scoreSig(15 downto 12),
			   Out0 => AhexU);	
HexA_L : HexDriver
	port map ( In0 => scoreSig(11 downto 8),
			   Out0 => AhexL);			
			   
HexB_U : HexDriver
	port map ( In0 => scoreSig(7 downto 4),
			   Out0 => BhexU);	
HexB_L : HexDriver
	port map ( In0 => scoreSig(3 downto 0),
			   Out0 => BhexL);					
			   	
		   
		   
	
Red <= redSig;
Blue <= blueSig;
Green <= greenSig;

vs <= vsSig;

end Behavioral;      
