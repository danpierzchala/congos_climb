library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

PACKAGE array_guySprite is
TYPE guySprite is array(26 downto 0, 26 downto 0) of integer;
END array_guySprite;
