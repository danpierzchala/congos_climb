library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

PACKAGE array_platPos is
TYPE platArray is array(0 to 7) of std_logic_vector(9 downto 0);
END array_platPos;

